`ifndef TB_PKG
`define TB_PKG
`include "uvm_macros.svh"
package tb_pkg;
    import uvm_pkg::*;
    `include "agent.sv"
    `include "env.sv"
    `include "test.sv"
endpackage
`endif
